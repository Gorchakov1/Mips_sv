`ifndef _MY_DEF
`define _MY_DEF

        `define OP_ADD		 4'b0001
	`define OP_MOV		 4'b0010
	`define OP_CMP		 4'b0011
	`define OP_SEE		 4'b0100
	`define OP_OR		  4'b0101
	`define OP_AND		 4'b0110
	`define OP_JMP   4'b0111
	`define OP_IN		  4'b1001
	`define OP_WR    4'b1010
	`define OP_JN    4'b1011
	`define OP_INC   4'b1100
	`define OP_DEC   4'b1101
	`define OP_END   4'b1110
        `define OP_JR    4'b1111	
`endif
	
